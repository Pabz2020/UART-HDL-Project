/*
 UART TX Controller
 Sends 1 byte of data serially: Start bit, 8 data bits (LSB first), Stop bit

 Inputs:
 - clk         : Baud rate clock tick (from baudRateGenerator)
 - reset_n     : Active-low asynchronous reset
 - i_Tx_Byte   : 8-bit data byte to send
 - i_Tx_Ready  : Signal to start transmission (pulse or held high)

 Outputs:
 - o_Tx_Data   : Serial UART TX output line
 - o_Tx_Done   : Pulses high for 1 clock tick after transmitting a byte
 - o_Tx_Active : High while transmission is in progress

*/

module uart_tx_controller(
    input        clk,
    input        reset_n,
    input  [7:0] i_Tx_Byte,
    input        i_Tx_Ready,
    output       o_Tx_Done,
    output       o_Tx_Active,
    output       o_Tx_Data
);

    // FSM states
    localparam UART_TX_IDLE  = 3'b000;
    localparam UART_TX_START = 3'b001;
    localparam UART_TX_DATA  = 3'b010;
    localparam UART_TX_STOP  = 3'b011;

    reg [2:0]  r_State      = UART_TX_IDLE;
    reg [2:0]  r_Bit_Index  = 0;
    reg        r_Tx_Data    = 1'b1;  // Idle line is logic HIGH
    reg        r_Tx_Done    = 1'b0;
    reg        r_Tx_Active  = 1'b0;

    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            r_State     <= UART_TX_IDLE;
            r_Bit_Index <= 3'd0;
            r_Tx_Data   <= 1'b1;
            r_Tx_Done   <= 1'b0;
            r_Tx_Active <= 1'b0;
        end else begin
            case (r_State)
                UART_TX_IDLE: begin
                    r_Tx_Done   <= 1'b0;
                    r_Tx_Data   <= 1'b1;  // Idle state line is HIGH
                    r_Bit_Index <= 3'd0;
                    r_Tx_Active <= 1'b0;
                    if (i_Tx_Ready) begin
                        r_State     <= UART_TX_START;
                        r_Tx_Active <= 1'b1;
                    end
                end

                UART_TX_START: begin
                    r_Tx_Data <= 1'b0;  // Start bit = 0
                    r_State   <= UART_TX_DATA;
                end

                UART_TX_DATA: begin
                    r_Tx_Data <= i_Tx_Byte[r_Bit_Index];
                    if (r_Bit_Index < 7) begin
                        r_Bit_Index <= r_Bit_Index + 1;
                    end else begin
                        r_Bit_Index <= 3'd0;
                        r_State     <= UART_TX_STOP;
                    end
                end

                UART_TX_STOP: begin
                    r_Tx_Data   <= 1'b1;  // Stop bit = 1
                    r_Tx_Done   <= 1'b1;  // Signal done for 1 clock
                    r_Tx_Active <= 1'b0;
                    r_State     <= UART_TX_IDLE;
                end

                default: begin
                    r_State <= UART_TX_IDLE;
                end
            endcase
        end
    end

    assign o_Tx_Data   = r_Tx_Data;
    assign o_Tx_Done   = r_Tx_Done;
    assign o_Tx_Active = r_Tx_Active;

endmodule
